`include "defines.svh"
module eth_port_fifo 
    (
        input clk,
        input rstn,
        input wr_en,
        input rd_en,
        input [`FIFO_WIDTH -1: 0] data_in,
        output reg [`FIFO_WIDTH -1: 0] data_out,
        output empty, full,
        output reg valid

    );

    reg [`FIFO_WIDTH -1: 0]mem[`FIFO_DEPTH -1: 0];
    bit [3:0] wr_ptr = 0;
    bit [3:0] rd_ptr = 0;

    bit empty_temp = 1'b1;
    bit full_temp = 1'b0;

    assign empty = empty_temp;
    assign full = full_temp;

    always @(*)
    begin
        if((wr_ptr == 0 && rd_ptr ==0) || (wr_ptr == rd_ptr))
            empty_temp = 1'b1;
        else 
            empty_temp = 1'b0;
        if(wr_ptr == `FIFO_DEPTH && rd_ptr ==0)
            full_temp = 1'b1;
        else
            full_temp = 1'b0;
    end

    always @(posedge clk)
    begin
        if(!rstn)
        begin
            data_out <= 'b0;
            wr_ptr <= 0;
            rd_ptr <= 0;
            valid <= 0;
            for(int i=0; i < `FIFO_DEPTH -1; i++)
            begin
                mem[i] <= 'b0;
            end
        end
        else
        begin
            if(wr_en)
            begin
                if(~full)
                begin
                    mem[wr_ptr] <= data_in;
                    $display("SW_DEBUG FIFO: data = %h filled in fifo loc %h \n",mem[wr_ptr], wr_ptr);
                    if(wr_ptr == `FIFO_DEPTH -1)
                    begin
                        $display("SW_DEBUG FIFO: wr_ptr reached the end of fifo");
                        wr_ptr <= 0;
                    end
                    else
                        wr_ptr <= wr_ptr +1;
                end
                else
                begin
                    $display("SW_DEBUG FIFO: FIFO is full \n");
                end
            end
            else if(rd_en)
            begin
                if(~empty)
                begin
                    data_out <= mem[rd_ptr];
                    valid <= 'b1;
                    if(rd_ptr == `FIFO_DEPTH -1)
                    begin
                        $display("SW_DEBUG FIFO: rd_ptr reached the end of fifo");
                        rd_ptr <= 0;
                    end
                    else
                        rd_ptr = rd_ptr +1;
                end
                else 
                begin
                    $display("SW_DEBUG FIFO: FIFO is empty \n");
                end
            end
        end
        if(valid == 1'b1)
            valid <= 1'b0;
    end

endmodule
