`define FIFO_DEPTH 10
`define FIFO_WIDTH 66
`define DATA_WIDTH 32
`define PORT_COUNT 2
